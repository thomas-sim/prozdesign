library ieee;
use ieee.std_logic_1164.all;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package from input file : seven_display.hex
-- ---------------------------------------------------------------------------------
package pkg_instrmem is

	type t_instrMem   is array(0 to 4096-1) of std_logic_vector(15 downto 0);
	constant PROGMEM : t_instrMem := (
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0010011111111111",
		"1110001111100011",
		"1000000100000000",
		"1110001111100110",
		"1000000100010000",
		"1110001111100101",
		"1000001100000000",
		"1110001111101000",
		"1000001100010000",
		"1100111111110111",
		
		others => (others => '0')
	);

end package pkg_instrmem;
