library ieee;
use ieee.std_logic_1164.all;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
package pkg_instrmem is

	type t_instrMem   is array(0 to 512-1) of std_logic_vector(15 downto 0);
	constant PROGMEM : t_instrMem := (
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"0000000000000000",
		"1110010100001010",
		"0010111000100000",
		"0010010000010001",
		"1110000000011000",
		"0000110000100010",
		"1111010000001000",
		"1001010000010011",
		"1001010100011010",
		"1111011111011001",
		"1100111111111111",
		
		others => (others => '0')
	);

end package pkg_instrmem;
